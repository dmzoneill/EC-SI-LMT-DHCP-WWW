IXA00366430 00:25:b3:ca:5b:96 10.243.18.216 /BLANK/ROOT/PATH
IXA00342559 00:22:64:33:59:37 10.243.18.123 /BLANK/ROOT/PATH
IXA00342560 00:23:7D:1B:AE:A6 10.243.18.131 /BLANK/ROOT/PATH
IXA00342561 00:23:7D:1B:B1:DC 10.243.18.137 /BLANK/ROOT/PATH
IXA00366508 00:09:6B:07:F0:FB 10.243.18.219 /BLANK/ROOT/PATH
IXA00384905 00:1e:67:2c:78:f7 10.243.18.63 /BLANK/ROOT/PATH
IXA00369888 00:E0:86:18:3A:A5 10.243.18.169 /BLANK/ROOT/PATH
IXA00369889 00:E0:86:17:00:32 10.243.18.221 /BLANK/ROOT/PATH
IXA00369890 00:e0:86:1b:bf:36 10.243.18.127 /BLANK/ROOT/PATH
IXA00369703 70:71:BC:DC:D0:1B 10.243.18.230 /BLANK/ROOT/PATH
IXA00368470 00:15:17:A1:C2:7F 10.243.18.89 /BLANK/ROOT/PATH
IXA00369309 78:2b:cb:af:1f:79 10.243.18.213 /BLANK/ROOT/PATH
IXA00378137 00:1E:67:3C:A3:7C 10.243.18.73 /BLANK/ROOT/PATH
IXA00370123 00:E0:86:18:26:58 10.243.18.117 /BLANK/ROOT/PATH
IXA00370127 00:E0:86:18:21:4E 10.243.18.205 /BLANK/ROOT/PATH
IXA00370137 00:E0:86:16:C4:2E 10.243.18.51 /BLANK/ROOT/PATH
IXA00370141 00:E0:86:18:3A:9A 10.243.18.180 /BLANK/ROOT/PATH
IXA00373698 00:1E:67:3C:77:8A 10.243.18.167 /BLANK/ROOT/PATH
IXA00386386 00:1E:67:43:3F:27 10.243.18.93 /BLANK/ROOT/PATH
IXA00384904 00:13:20:fd:f9:3d 10.243.18.113 /BLANK/ROOT/PATH
IXA00370130 00:E0:86:18:3A:9F 10.243.18.129 /BLANK/ROOT/PATH
IXA00370367 18:03:73:C8:48:10 10.243.18.223 /BLANK/ROOT/PATH
IXA00371268 18:03:73:D9:71:D1 10.243.18.162 /BLANK/ROOT/PATH
IXA00368859 00:01:80:7C:C6:7D 10.243.18.151 /BLANK/ROOT/PATH
IXA00370133 00:E0:86:16:C4:36 10.243.18.248 /BLANK/ROOT/PATH
IXA00370385 00:E0:86:18:3B:78 10.243.18.159 /BLANK/ROOT/PATH
IXA00370839 E0:69:95:EB:75:CD 10.243.18.233 /BLANK/ROOT/PATH
IXA00379666 00:1E:67:43:4A:3A 10.243.18.106 /BLANK/ROOT/PATH
IXA00385949 00:1E:67:59:77:AB 10.243.18.28 /BLANK/ROOT/PATH
IXA00380745 00:1B:21:00:6C:45 10.243.18.157 /BLANK/ROOT/PATH
IXA00379576 E0:69:95:D3:0D:1B 10.243.18.103 /BLANK/ROOT/PATH
IXA00379771 00:e0:86:1b:bf:33 10.243.18.243 /BLANK/ROOT/PATH
IXA00370365 18:03:73:C6:EE:F1 10.243.18.165 /BLANK/ROOT/PATH
IXA00371766 00:1E:67:2C:75:82 10.243.18.182 /BLANK/ROOT/PATH
IXA00379582 00:11:22:33:44:55 10.243.18.178 /BLANK/ROOT/PATH
IXA00384834 00:13:20:FF:1C:E2 10.243.18.246 /BLANK/ROOT/PATH
IXA00379955 00:1e:67:43:40:0E 10.243.18.130 /BLANK/ROOT/PATH
IXA00379496 00:1e:67:43:48:65 10.243.18.235 /BLANK/ROOT/PATH
IXA00370364 00:1b:21:8c:73:f0 10.243.18.164 /BLANK/ROOT/PATH
IXA00372153 E0:69:95:D3:05:47 10.243.18.87 /BLANK/ROOT/PATH
IXA00372516 38:60:77:12:74:C0 10.243.18.254 /BLANK/ROOT/PATH
IXA00380742 68:05:ca:08:6b:e4 10.243.18.202 /BLANK/ROOT/PATH
IXA00382993 00:1E:67:59:81:A8 10.243.18.100 /BLANK/ROOT/PATH
IXA00371572 00:1e:67:2c:77:9e 10.243.18.97 /BLANK/ROOT/PATH
IXA00384488 78:2B:CB:94:F8:E7 10.243.18.66 /BLANK/ROOT/PATH
IXA00384443 00:1E:67:43:44:59 10.243.18.143 /BLANK/ROOT/PATH
IXA00384442 9C:8E:99:52:63:DE 10.243.18.181 /BLANK/ROOT/PATH
IXA00384441 00:1E:67:3C:76:21 10.243.18.251 /BLANK/ROOT/PATH
IXA00365684 00:15:17:be:28:5e 10.243.18.135 /BLANK/ROOT/PATH
IXA00370838 E0:69:95:E4:F6:D2 10.243.18.161 /BLANK/ROOT/PATH
IXA00386010 00:1e:67:59:81:a9 10.243.18.215 /BLANK/ROOT/PATH
IXA00380551 90:2B:34:5B:1B:E6 10.243.18.14 /BLANK/ROOT/PATH
IXA00386024 78:54:2E:E6:0A:E9 10.243.18.163 /BLANK/ROOT/PATH
IXA00386025 00:13:20:fd:df:55 10.243.18.146 /BLANK/ROOT/PATH
IXA00386030 e0:db:55:b9:5d:ac 10.243.18.252 /BLANK/ROOT/PATH
IXA00380743 00:15:17:BE:26:DB 10.243.18.134 /BLANK/ROOT/PATH
IXA00384452 00:1e:67:59:78:30 10.243.18.119 /BLANK/ROOT/PATH
IXA00384465 00:1B:21:1B:FD:A6 10.243.18.152 /BLANK/ROOT/PATH
IXA00368862 00:01:80:7C:9E:CD 10.243.18.53 /BLANK/ROOT/PATH
IXA00384535 94:DE:80:6E:F5:89 10.243.18.199 /BLANK/ROOT/PATH
IXA00384536 94:DE:80:6D:04:3A 10.243.18.201 /BLANK/ROOT/PATH
IXA00382993 00:1E:67:59:81:A8 10.243.18.6 /BLANK/ROOT/PATH
IXA00367097 00:15:17:EA:C1:05 10.243.18.7 /BLANK/ROOT/PATH
IXA00384508 00:1E:67:3C:79:82 10.243.18.217 /BLANK/ROOT/PATH
IXA00371415 00:1E:67:2C:77:C7 10.243.18.249 /BLANK/ROOT/PATH
IXA00384907 00:15:17:af:76:68 10.243.18.214 /BLANK/ROOT/PATH
IXA00384908 78:ac:c0:be:4a:45 10.243.18.191 /BLANK/ROOT/PATH
IXA00384906 18:03:73:c6:bc:d6 10.243.18.239 /BLANK/ROOT/PATH
IXA00372535 E0:69:95:EB:3D:06 10.243.18.118 /BLANK/ROOT/PATH
IXA00372465 E0:69:95:EB:48:2E 10.243.18.140 /BLANK/ROOT/PATH
IXA00380360 00:22:4d:80:f4:06 10.243.18.156 /BLANK/ROOT/PATH
IXA00383020 00:13:20:FD:23:03 10.243.18.225 /BLANK/ROOT/PATH
IXA00373699 00:1E:67:3C:77:9F 10.243.18.172 /BLANK/ROOT/PATH
IXA00384451 00:1C:C4:73:C7:70 10.243.18.174 /BLANK/ROOT/PATH
IXA00379736 00:1e:67:49:B0:CA 10.243.18.176 /BLANK/ROOT/PATH
IXA00386352 00:1E:67:43:46:B3 10.243.18.253 /BLANK/ROOT/PATH
IXA00384578 00:08:A2:09:04:19 10.243.18.23 /BLANK/ROOT/PATH
IXA00385264 1c:6f:65:9c:fa:a1 10.243.18.196 /BLANK/ROOT/PATH
IXA00369304 78:2B:CB:AF:1E:C1 10.243.18.5 /BLANK/ROOT/PATH
IXA00379448 00:1E:67:43:46:AD 10.243.18.19 /BLANK/ROOT/PATH
IXA00384024 00:E0:86:1B:BF:3B 10.243.18.155 /BLANK/ROOT/PATH
IXA00384434 18:03:73:D9:70:AC 10.243.18.179 /BLANK/ROOT/PATH
IXA00384878 00:1E:67:3c:79:43 10.243.18.244 /BLANK/ROOT/PATH
IXA00378942 00:1E:67:43:48:96 10.243.18.108 /BLANK/ROOT/PATH
IXA00386175 00:1E:67:59:77:19 10.243.18.195 /BLANK/ROOT/PATH
IXA00384880 00:1B:21:43:51:34 10.243.18.184 /BLANK/ROOT/PATH
IXA00378943 00:1E:67:3C:A3:0D 10.243.18.231 /BLANK/ROOT/PATH
